module adder_4(pc, new_pc);
	new_pc = pc + 4;
endmodule